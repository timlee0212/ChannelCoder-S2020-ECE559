`timescale 1ns/1ps
module tb_full();
//Input Ports
reg clk, reset, tb_in, wreq_tb, wreq_size;

reg[15:0] tb_size_in;

//Output Ports
wire ck_out, zk_out, zk_prime_out;

coder_stack_top test_obj(
	.clk(clk),
	.reset(reset), 
	.tb_in(tb_in), 
	.wreq_data(wreq_tb), 
	.tb_size_in(tb_size_in), 
	.wreq_size(wreq_size),
	.xk_out(xk_out), 
	.zk_out(zk_out), 
	.zk_prime_out(zk_prime_out)
);


integer length = 7010;
integer iterations = 7250, i, k;

wire[7009:0] input_vector = 7010'b01010111010000111110001010010101011011111101101010101110000010110010001010010000111111001100011100010000100001101111000100101011010111100000011001011101100101101111101010011010111110011011000111011110010111000101101111001000111101001001101100111001000001111101001000000001000101001101101001001100000100111010000101110001100011011000111100010101101111111110110011100010111000101110001001110010101111010110100011000101010011011000001010011011001111110110011101100000111000111011111110100000011000100001001001001111011000010000101101010000010001110100011000111001100100001011000101010101000010101001101001001101011000010111010010011110010000010110010100010001111011000001010100100110100000100110011011011000111100111110000000000000110011001101001010101001001000100000101011110100100101111110100110001101000011011011000001001011100100101100001001101001101111100000010010111000010100000101010100011100111111101011111001011111110101110010110010101011010001110000001011111110100111011101011100000000011000111101010110111110000110010010001111000111110100010110010101111000000001000010001111101101010010011001100011000110111111111100110001011101100101101011111101001010110001101000101111110110011001000010000011011101101101100010111001101011100110010100001010111000000110011011110000100100100100011111011011100111000000011100000101010001000000001011001000000110111111001110011010000000101111011111010000010101110011111010101010110000110010101100000110101000100010110001110001110010001100011100011101100101100111001001110011001110000100011001001001010101110011101100000101000000100000100100111010010001110010011110000000101101100001010000011011001111010111001010001110111101000110101000011100000011111111010111010001111100001101101100101100101100010100011110101110010111000100100100100100111100001101011000100011011010001100010101101011000001111100010000000100100011011001101101111010111111110010000010111101001111001111101101111101001010011110001110110010110000011111110011100101111101111101101011011100000101100100101100011100011100101100101011110011001111001011000011011110100101110011010100111101111100000111111100101101101000101001111100101001000011010111011101010010011100001101110101111101111110001111000110000000110011001001110000011100010000110000111110110001010101001110111111000101111111110001010101001010101111011101011110011110101101000100000111011001011010010111111001100100101000001000011111111110110111000110000101110111010101100101001011001110001001011010001000111100101101101000111001001111111100011000010000111001010100110011000101010001011110110101101001011001110010011001001000001001100010100001010001011000000011001001000011010010010101110100100011011010001011001011001000111000000111100110100111010100011100000000110111110101110010110000111010101111000100110110010101101001000100001010110100111000001110011001111010011100101111110001010111000010101101011100001001001110010000101111001100110010010001110110111110010010111111011110101001110101010100110100101010110010001101010111111111100001110111010011001011100000000100000111000100100101011000000101001000000011101011100001010010101010100001000101011100000010111011110110010100000100000100011111101101100001111001011011100011100000000111111101100000010111110101101011111011101111100111011110000101111111100000011111100110101010100000000000100100000110011101001001100100010001001101101111101110000111101000111001011011111010101010101110011000010000110011101100011010011011010010010001100001100110010011100001000010000100001010110000110101101110001011100101010010001110001011100100000101000010101011100111101111011000111010111000011110100101010001001101011010010010100100011100110001011110110010101011011011001010011111110011011100001111010001100010100011000000101011111101100101101011110100001010010001010011000000111001010101010101011100111101001011111000111101000110100101000101100010101110001000100000111101001010101110011010000001010000110111001010000001010100110001001001101111000000010100100101101110001100010010101111001010101010100101000000110101111001111101111011000101110100101101100010001100110011001111111011111001010101100110011111101001010001110001101101000101011111000111101100110101001000101010101001010000100011001110011000001111110100010011001101111011011001101100111011001001010011001010001011001101101010010000010001010010000100000001100011101101101110000010010011001101011101011000100111100101001111010010110111101100110011011100011001110101110101011110101000010111111001101000000100110001111001111101110001010000100100100100000110001100000011100111100011110110111001110101000111101001100011111001111110011000100101000000010101001010001111101101000011011111110000000001110111111001010111100100011111101000010100000101010110101000010110111101110000111111100110011110110000100111101100100101001111100001110000100001110011000000000011110100001001100011011111110100101100101010000101101001101101100111010000000100011110010000110011010010000110110010100010111001010011111011111100110001011101111111100001110111001100100001101000111110001110000000111100011111000001001111111111110010111001000011101101100000010101000110011000011110110000111111101100100001110010011000000001100010001100000110010111010110111011011000101001010000011001111001100011111100100100011000001010001001110001000001100001000110010110100010100111111010101111111110100010110100111100011111111011011101010000010110010010000111101111001111010101010101101110011011000111011101100010101101011011100000000000101011011000111000010100110000101101011101000110101101100000001000001000011011110110110000000111101010010110101101101110000110010100111100000001001001101001000000100011101000100101011000010101001010011011101011000110111000101111011001000010010111111001011001101110000101000000010101000000101000010001111111100000100001111101000010000110001101100110010000000100010011001111010011011100001000010110010100001101110101001100010110001111001111111110001110011011010011001111100100111000010000111110010101111000101101000001010100111111101000110000011110011011001011011001001110100100101100010000001101011110100000101100001100101000100100100010110000001110011000010000011010101011110110100010101111001110110111101101111100000100010001111111110000000100011000011110101111111000011000111101110100111000011000110101001100110011110001001010001110000111001100101010110000110110000000000000101001001000111111111100010000101111000001110001000100101101000001011100110101101001010110110001111110001110110110000100011010100010100100010111111110011000010000100011100011111101011110110111011011101011110000101011001111111110010001000101000000100000100001000010111100100101001110110110100111000111001000000110110100010010110010011110101110001111000010000101100101011011100011100010011001101111100011100111001001111001100000011001001100100101011100000000110100011001001010111101010101111001111011011111001001110001001011111100010000010111010001010010011001011011010101001001001001000000010010101110110011010101111000100100100000000100000111010100101011010111100010010111001111101110;

//Clock Generator
initial clk=1'b0;
always #5 clk=~clk;

//Power-on Reset
initial
begin
		reset = 1'b1;
#20 	reset = 1'b0;
end


initial
begin	
	wreq_size = 1'b0;
	wreq_tb = 1'b0;
	tb_size_in = 16'h0;
	tb_in = 1'b0;
end

initial
begin
#50	wreq_size = 1'b1;
		tb_size_in = length;
#15	wreq_size = 1'b0;
#25	wreq_tb = 1'b1;
#5
	i = 0;
	k = -1;
	while (i < iterations)
	begin
		//#10 
		
		if (i < 7010) 
			tb_in = input_vector[i];
		else
			tb_in = 0;
		#10 i = i + 1;
	end
	wreq_tb = 1'b0;
end
endmodule
