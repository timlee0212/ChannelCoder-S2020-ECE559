`timescale 1ns/1ps
module tb_full();
//Input Ports
reg clk, reset, wreq_tb, wreq_size;
reg[7:0] tb_in;

reg[11:0] tb_size_in;

//Output Ports
wire[7:0] xk_out, zk_out, zk_prime_out, d_cbs_out;
wire out_valid;

coder_stack_top test_obj(
	.clk(clk),
	.reset(reset), 
	.tb_in(tb_in), 
	.wreq_data(wreq_tb), 
	.tb_size_in(tb_size_in), 
	.wreq_size(wreq_size),
	.xk_out(xk_out), 
	.zk_out(zk_out), 
	.zk_prime_out(zk_prime_out),
	.out_valid(out_valid)
);


integer length = 878;
integer iterations = 925, i, k;


integer f_xk, f_zk, f_zk_p;

initial begin
	f_xk = $fopen("xk.txt", "w");
	f_zk = $fopen("zk.txt", "w");
	f_zk_p = $fopen("zk_p.txt", "w");
end


wire[7023:0] input_vector = 7024'b0101011101000011111000101001010101101111110110101010111000001011001000101001000011111100110001110001000010000110111100010010101101011110000001100101110110010110111110101001101011111001101100011101111001011100010110111100100011110100100110110011100100000111110100100000000100010100110110100100110000010011101000010111000110001101100011110001010110111111111011001110001011100010111000100111001010111101011010001100010101001101100000101001101100111111011001110110000011100011101111111010000001100010000100100100111101100001000010110101000001000111010001100011100110010000101100010101010100001010100110100100110101100001011101001001111001000001011001010001000111101100000101010010011010000010011001101101100011110011111000000000000011001100110100101010100100100010000010101111010010010111111010011000110100001101101100000100101110010010110000100110100110111110000001001011100001010000010101010001110011111110101111100101111111010111001011001010101101000111000000101111111010011101110101110000000001100011110101011011111000011001001000111100011111010001011001010111100000000100001000111110110101001001100110001100011011111111110011000101110110010110101111110100101011000110100010111111011001100100001000001101110110110110001011100110101110011001010000101011100000011001101111000010010010010001111101101110011100000001110000010101000100000000101100100000011011111100111001101000000010111101111101000001010111001111101010101011000011001010110000011010100010001011000111000111001000110001110001110110010110011100100111001100111000010001100100100101010111001110110000010100000010000010010011101001000111001001111000000010110110000101000001101100111101011100101000111011110100011010100001110000001111111101011101000111110000110110110010110010110001010001111010111001011100010010010010010011110000110101100010001101101000110001010110101100000111110001000000010010001101100110110111101011111111001000001011110100111100111110110111110100101001111000111011001011000001111111001110010111110111110110101101110000010110010010110001110001110010110010101111001100111100101100001101111010010111001101010011110111110000011111110010110110100010100111110010100100001101011101110101001001110000110111010111110111111000111100011000000011001100100111000001110001000011000011111011000101010100111011111100010111111111000101010100101010111101110101111001111010110100010000011101100101101001011111100110010010100000100001111111111011011100011000010111011101010110010100101100111000100101101000100011110010110110100011100100111111110001100001000011100101010011001100010101000101111011010110100101100111001001100100100000100110001010000101000101100000001100100100001101001001010111010010001101101000101100101100100011100000011110011010011101010001110000000011011111010111001011000011101010111100010011011001010110100100010000101011010011100000111001100111101001110010111111000101011100001010110101110000100100111001000010111100110011001001000111011011111001001011111101111010100111010101010011010010101011001000110101011111111110000111011101001100101110000000010000011100010010010101100000010100100000001110101110000101001010101010000100010101110000001011101111011001010000010000010001111110110110000111100101101110001110000000011111110110000001011111010110101111101110111110011101111000010111111110000001111110011010101010000000000010010000011001110100100110010001000100110110111110111000011110100011100101101111101010101010111001100001000011001110110001101001101101001001000110000110011001001110000100001000010000101011000011010110111000101110010101001000111000101110010000010100001010101110011110111101100011101011100001111010010101000100110101101001001010010001110011000101111011001010101101101100101001111111001101110000111101000110001010001100000010101111110110010110101111010000101001000101001100000011100101010101010101110011110100101111100011110100011010010100010110001010111000100010000011110100101010111001101000000101000011011100101000000101010011000100100110111100000001010010010110111000110001001010111100101010101010010100000011010111100111110111101100010111010010110110001000110011001100111111101111100101010110011001111110100101000111000110110100010101111100011110110011010100100010101010100101000010001100111001100000111111010001001100110111101101100110110011101100100101001100101000101100110110101001000001000101001000010000000110001110110110111000001001001100110101110101100010011110010100111101001011011110110011001101110001100111010111010101111010100001011111100110100000010011000111100111110111000101000010010010010000011000110000001110011110001111011011100111010100011110100110001111100111111001100010010100000001010100101000111110110100001101111111000000000111011111100101011110010001111110100001010000010101011010100001011011110111000011111110011001111011000010011110110010010100111110000111000010000111001100000000001111010000100110001101111111010010110010101000010110100110110110011101000000010001111001000011001101001000011011001010001011100101001111101111110011000101110111111110000111011100110010000110100011111000111000000011110001111100000100111111111111001011100100001110110110000001010100011001100001111011000011111110110010000111001001100000000110001000110000011001011101011011101101100010100101000001100111100110001111110010010001100000101000100111000100000110000100011001011010001010011111101010111111111010001011010011110001111111101101110101000001011001001000011110111100111101010101010110111001101100011101110110001010110101101110000000000010101101100011100001010011000010110101110100011010110110000000100000100001101111011011000000011110101001011010110110111000011001010011110000000100100110100100000010001110100010010101100001010100101001101110101100011011100010111101100100001001011111100101100110111000010100000001010100000010100001000111111110000010000111110100001000011000110110011001000000010001001100111101001101110000100001011001010000110111010100110001011000111100111111111000111001101101001100111110010011100001000011111001010111100010110100000101010011111110100011000001111001101100101101100100111010010010110001000000110101111010000010110000110010100010010010001011000000111001100001000001101010101111011010001010111100111011011110110111110000010001000111111111000000010001100001111010111111100001100011110111010011100001100011010100110011001111000100101000111000011100110010101011000011011000000000000010100100100011111111110001000010111100000111000100010010110100000101110011010110100101011011000111111000111011011000010001101010001010010001011111111001100001000010001110001111110101111011011101101110101111000010101100111111111001000100010100000010000010000100001011110010010100111011011010011100011100100000011011010001001011001001111010111000111100001000010110010101101110001110001001100110111110001110011100100111100110000001100100110010010101110000000011010001100100101011110101010111100111101101111100100111000100101111110001000001011101000101001001100101101101010100100100100100000001001010111011001101010111100010010010000000010000011101010010101101011110001001011100111110111001110000111100;

//Clock Generator
initial clk=1'b0;
always #5 clk=~clk;


reg prev_out_valid;
always @(posedge clk) begin
	if (out_valid) begin
		$fwrite(f_xk, "%8b\n", xk_out);
		$fwrite(f_zk, "%8b\n", zk_out);
		$fwrite(f_zk_p, "%8b\n", zk_prime_out);
		prev_out_valid = out_valid;
	end
	else begin
		if (prev_out_valid) begin
			$fclose(f_xk);
			$fclose(f_zk);
			$fclose(f_zk_p);
			$stop();
		end
	end
end


//Power-on Reset
initial
begin
		reset = 1'b1;
#20 	reset = 1'b0;
end


initial
begin	
	wreq_size = 1'b0;
	wreq_tb = 1'b0;
	tb_size_in = 16'h0;
	tb_in = 1'b0;
end

initial
begin
#50	wreq_size = 1'b1;
		tb_size_in = length;
#15	wreq_size = 1'b0;
#25	wreq_tb = 1'b1;
#5
	i = 0;
	k = -1;
	while (i < iterations)
	begin
		//#10 
		
		if (i < length) 
			tb_in = input_vector[i * 8 +: 8];
		else
			tb_in = 0;
		#10 i = i + 1;
	end
	wreq_tb = 1'b0;
end
endmodule
